.SUBCKT NAND3 A B C OUT VDD VSS
MM0 OUT A VDD VDD p_18 W=2u L=180.00n
MM1 OUT B VDD VDD p_18 W=2u L=180.00n
MM2 OUT C VDD VDD p_18 W=2u L=180.00n
MM3 OUT C net1 VSS n_18 W=3u L=180.00n
MM4 net1 B net0 VSS n_18 W=3u L=180.00n
MM5 net0 A VSS VSS n_18 W=3u L=180.00n
.ENDS

.SUBCKT NOR2 A B OUT VDD VSS
MM0 net0 A VDD VDD p_18 W=40u L=180.00n
MM1 OUT B net0 VDD p_18 W=40u L=180.00n
MM2 OUT B VSS VSS n_18 W=10u L=180.00n
MM3 OUT A VSS VSS n_18 W=10u L=180.00n
.ENDS


.SUBCKT B IN OUT VDD VSS
X1 VDD VDD VDD net0 VDD VSS NAND3
X2 IN VDD VDD net1 VDD VSS NAND3
X3 net1 net0 OUT VDD VSS NOR2
.ENDS
