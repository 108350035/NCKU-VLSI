.SUBCKT INV IN OUT VDD VSS
MM0 OUT IN VDD VDD p_18 W=6u L=180.00n
MM1 OUT IN VSS VSS n_18 W=2u L=180.00n
.ENDS

.SUBCKT INV_CHAIN pulse_in pulse_out VDD VSS
X1 pulse_in A VDD VSS INV
X2 A IN VDD VSS INV M=M1
X3 IN OUT VDD VSS INV M=M2
X4 OUT B VDD VSS INV M=M3
X5 B pulse_out VDD VSS INV M=M4
.ENDS


