* File: ring_osc.pex.spi
* Created: Tue Apr 15 12:12:30 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "ring_osc.pex.spi.pex"
.subckt ring_osc  IN VSS VDD
* 
* VDD	VDD
* VSS	VSS
* IN	IN
mx1.MM4 N_NET0_x1.MM4_d N_IN_x1.MM4_g N_VSS_x1.MM4_s N_VSS_x1.MM4_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx1.MM4@2 N_NET0_x1.MM4@2_d N_IN_x1.MM4@2_g N_VSS_x1.MM4@2_s N_VSS_x1.MM4_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx2.MM4 N_NET1_x2.MM4_d N_NET0_x2.MM4_g N_VSS_x2.MM4_s N_VSS_x1.MM4_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx2.MM4@2 N_NET1_x2.MM4@2_d N_NET0_x2.MM4@2_g N_VSS_x2.MM4@2_s N_VSS_x1.MM4_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx3.MM4 N_NET2_x3.MM4_d N_NET1_x3.MM4_g N_VSS_x3.MM4_s N_VSS_x1.MM4_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx3.MM4@2 N_NET2_x3.MM4@2_d N_NET1_x3.MM4@2_g N_VSS_x3.MM4@2_s N_VSS_x1.MM4_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx4.MM4 N_NET3_x4.MM4_d N_NET2_x4.MM4_g N_VSS_x4.MM4_s N_VSS_x1.MM4_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx4.MM4@2 N_NET3_x4.MM4@2_d N_NET2_x4.MM4@2_g N_VSS_x4.MM4@2_s N_VSS_x1.MM4_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx5.MM4 N_IN_x5.MM4_d N_NET3_x5.MM4_g N_VSS_x5.MM4_s N_VSS_x1.MM4_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx5.MM4@2 N_IN_x5.MM4@2_d N_NET3_x5.MM4@2_g N_VSS_x5.MM4@2_s N_VSS_x1.MM4_b N_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mx1.MM0 N_NET0_x1.MM0_d N_IN_x1.MM0_g N_VDD_x1.MM0_s N_VDD_x1.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx1.MM0@2 N_NET0_x1.MM0@2_d N_IN_x1.MM0@2_g N_VDD_x1.MM0@2_s N_VDD_x1.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx2.MM0 N_NET1_x2.MM0_d N_NET0_x2.MM0_g N_VDD_x2.MM0_s N_VDD_x1.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx2.MM0@2 N_NET1_x2.MM0@2_d N_NET0_x2.MM0@2_g N_VDD_x2.MM0@2_s N_VDD_x1.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx3.MM0 N_NET2_x3.MM0_d N_NET1_x3.MM0_g N_VDD_x3.MM0_s N_VDD_x1.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx3.MM0@2 N_NET2_x3.MM0@2_d N_NET1_x3.MM0@2_g N_VDD_x3.MM0@2_s N_VDD_x1.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx4.MM0 N_NET3_x4.MM0_d N_NET2_x4.MM0_g N_VDD_x4.MM0_s N_VDD_x1.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx4.MM0@2 N_NET3_x4.MM0@2_d N_NET2_x4.MM0@2_g N_VDD_x4.MM0@2_s N_VDD_x1.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx5.MM0 N_IN_x5.MM0_d N_NET3_x5.MM0_g N_VDD_x5.MM0_s N_VDD_x1.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mx5.MM0@2 N_IN_x5.MM0@2_d N_NET3_x5.MM0@2_g N_VDD_x5.MM0@2_s N_VDD_x1.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
*
.include "ring_osc.pex.spi.RING_OSC.pxi"
*
.ends
*
*
