.SUBCKT A3 A B C D E OUT VDD VSS
MM0 net0 B VSS VSS n_18 W=1u L=180.00n
MM1 net0 C VSS VSS n_18 W=1u L=180.00n
MM2 net0 D VSS VSS n_18 W=1u L=180.00n
MM3 net0 E VSS VSS n_18 W=1u L=180.00n
MM4 OUT A net0 VSS n_18 W=1u L=180.00n

MM5 OUT A VDD VDD p_18 W=3u L=180.00n
MM6 OUT B net1 VDD p_18 W=12u L=180.00n
MM7 net1 C net2 VDD p_18 W=12u L=180.00n
MM8 net2 D net3 VDD p_18 W=12u L=180.00n
MM9 net3 E VDD VDD p_18 W=12u L=180.00n
.ENDS

