* File: AND6_pseudo.pex.spi
* Created: Tue Apr 22 09:22:13 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "AND6_pseudo.pex.spi.pex"
.subckt nand6  VSS B A D C F E VDD OUT
* 
* OUT	OUT
* VDD	VDD
* E	E
* F	F
* C	C
* D	D
* A	A
* B	B
* VSS	VSS
MM1 N_NET1_MM1_d N_B_MM1_g N_NET0_MM1_s N_VSS_MM1_b N_18 L=1.8e-07 W=2.7e-06
+ AD=1.323e-12 AS=6.885e-13 PD=3.68e-06 PS=5.1e-07
MM2 N_NET0_MM2_d N_A_MM2_g N_VSS_MM2_s N_VSS_MM1_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.885e-13 AS=1.323e-12 PD=5.1e-07 PS=3.68e-06
MM4 N_NET3_MM4_d N_D_MM4_g N_NET2_MM4_s N_VSS_MM1_b N_18 L=1.8e-07 W=2.7e-06
+ AD=1.323e-12 AS=6.885e-13 PD=3.68e-06 PS=5.1e-07
MM5 N_NET2_MM5_d N_C_MM5_g N_VSS_MM5_s N_VSS_MM1_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.885e-13 AS=1.323e-12 PD=5.1e-07 PS=3.68e-06
MM7 N_NET5_MM7_d N_F_MM7_g N_NET4_MM7_s N_VSS_MM1_b N_18 L=1.8e-07 W=2.7e-06
+ AD=1.323e-12 AS=6.885e-13 PD=3.68e-06 PS=5.1e-07
MM8 N_NET4_MM8_d N_E_MM8_g N_VSS_MM8_s N_VSS_MM1_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.885e-13 AS=1.323e-12 PD=5.1e-07 PS=3.68e-06
MM12 N_OUT_MM12_d N_NET5_MM12_g N_VSS_MM12_s N_VSS_MM1_b N_18 L=1.8e-07
+ W=2.1e-06 AD=5.355e-13 AS=1.029e-12 PD=5.1e-07 PS=3.08e-06
MM12@2 N_OUT_MM12@2_d N_NET5_MM12@2_g N_VSS_MM12@2_s N_VSS_MM1_b N_18 L=1.8e-07
+ W=2.1e-06 AD=5.355e-13 AS=5.355e-13 PD=5.1e-07 PS=5.1e-07
MM11 N_OUT_MM11_d N_NET3_MM11_g N_VSS_MM11_s N_VSS_MM1_b N_18 L=1.8e-07
+ W=2.1e-06 AD=5.355e-13 AS=5.355e-13 PD=5.1e-07 PS=5.1e-07
MM11@2 N_OUT_MM11@2_d N_NET3_MM11@2_g N_VSS_MM11@2_s N_VSS_MM1_b N_18 L=1.8e-07
+ W=2.1e-06 AD=5.355e-13 AS=5.355e-13 PD=5.1e-07 PS=5.1e-07
MM10 N_OUT_MM10_d N_NET1_MM10_g N_VSS_MM10_s N_VSS_MM1_b N_18 L=1.8e-07
+ W=2.1e-06 AD=5.355e-13 AS=5.355e-13 PD=5.1e-07 PS=5.1e-07
MM10@2 N_OUT_MM10@2_d N_NET1_MM10@2_g N_VSS_MM10@2_s N_VSS_MM1_b N_18 L=1.8e-07
+ W=2.1e-06 AD=5.355e-13 AS=1.029e-12 PD=5.1e-07 PS=3.08e-06
MM0 N_NET1_MM0_d N_VSS_MM0_g N_VDD_MM0_s N_VDD_MM0_b P_18 L=1.8e-07 W=6.8e-07
+ AD=3.332e-13 AS=3.332e-13 PD=1.66e-06 PS=1.66e-06
MM3 N_NET3_MM3_d N_VSS_MM3_g N_VDD_MM3_s N_VDD_MM0_b P_18 L=1.8e-07 W=6.8e-07
+ AD=3.332e-13 AS=3.332e-13 PD=1.66e-06 PS=1.66e-06
MM6 N_NET5_MM6_d N_VSS_MM6_g N_VDD_MM6_s N_VDD_MM0_b P_18 L=1.8e-07 W=6.8e-07
+ AD=3.332e-13 AS=3.332e-13 PD=1.66e-06 PS=1.66e-06
MM9 N_OUT_MM9_d N_VSS_MM9_g N_VDD_MM9_s N_VDD_MM0_b P_18 L=1.8e-07 W=2.1e-06
+ AD=1.029e-12 AS=1.029e-12 PD=3.08e-06 PS=3.08e-06
*
.include "AND6_pseudo.pex.spi.AND6_PSEUDO.pxi"
*
.ends
*
*
