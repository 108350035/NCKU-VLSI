.SUBCKT NAND2 A B OUT VDD VSS
MM0 OUT A VDD VDD p_18 W=2.5u L=180.00n
MM1 OUT B VDD VDD p_18 W=2.5u L=180.00n
MM4 OUT B net0 VSS n_18 W=2.5u L=180.00n
MM5 net0 A VSS VSS n_18 W=2.5u L=180.00n
.ENDS

.SUBCKT NOR3 A B C OUT VDD VSS
MM0 net0 A VDD VDD p_18 W=56.98u L=180.00n
MM1 net1 B net0 VDD p_18 W=56.98u L=180.00n
MM2 OUT C net1 VDD p_18 W=56.98u L=180.00n
MM3 OUT C VSS VSS n_18 W=9.5u L=180.00n
MM4 OUT B VSS VSS n_18 W=9.5u L=180.00n
MM5 OUT A VSS VSS n_18 W=9.5u L=180.00n
.ENDS


.SUBCKT C IN OUT VDD VSS
X1 VDD VDD net0 VDD VSS NAND2
X2 VDD VDD net1 VDD VSS NAND2
X3 IN VDD net2 VDD VSS NAND2
X4 net2 net1 net0 OUT VDD VSS NOR3
.ENDS
