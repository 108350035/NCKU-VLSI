.SUBCKT INV IN OUT VDD VSS
MM0 OUT IN VDD VDD p_18 W=3u L=180.00n
MM4 OUT IN VSS VSS n_18 W=0.94u L=180.00n
.ENDS

.SUBCKT ring_osc IN VDD VSS
x1 IN net0 VDD VSS INV
x2 net0 net1 VDD VSS INV
x3 net1 net2 VDD VSS INV
x4 net2 net3 VDD VSS INV
x5 net3 IN VDD VSS INV
.ENDS

