*ttt
.SUBCKT NMOS D G S B
MM0 D G S B n_18 W=6u L=180.00n
.ENDS

.SUBCKT PMOS D G S B
MM0 D G S B p_18 W=15u L=180.00n
.ENDS
