************************************************************************
* auCdl Netlist:
* 
* Library Name:  mylib
* Top Cell Name: decoder
* View Name:     schematic
* Netlisted on:  Apr  6 22:54:44 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: mylib
* Cell Name:    decoder
* View Name:    schematic
************************************************************************

.SUBCKT decoder A B C D O1 O2 O3 O4 O5 O6 O7 O8 VDD VSS
*.PININFO A:I B:I C:I D:I VDD:I VSS:I O1:O O2:O O3:O O4:O O5:O O6:O O7:O O8:O
MM77 O1 net0143 VDD VDD p_18 W=1u L=180.00n
MM75 net0143 A VDD VDD p_18 W=1u L=180.00n
MM71 net0143 D VDD VDD p_18 W=1u L=180.00n
MM70 net0143 C VDD VDD p_18 W=1u L=180.00n
MM69 net0143 B VDD VDD p_18 W=1u L=180.00n
MM68 O2 net0145 VDD VDD p_18 W=1u L=180.00n
MM66 net0145 A VDD VDD p_18 W=1u L=180.00n
MM62 net0145 ~D VDD VDD p_18 W=1u L=180.00n
MM61 net0145 C VDD VDD p_18 W=1u L=180.00n
MM60 net0145 B VDD VDD p_18 W=1u L=180.00n
MM59 O3 net0107 VDD VDD p_18 W=1u L=180.00n
MM57 net0107 A VDD VDD p_18 W=1u L=180.00n
MM53 net0107 D VDD VDD p_18 W=1u L=180.00n
MM52 net0107 ~C VDD VDD p_18 W=1u L=180.00n
MM51 net0107 B VDD VDD p_18 W=1u L=180.00n
MM50 O4 net0109 VDD VDD p_18 W=1u L=180.00n
MM48 net0109 A VDD VDD p_18 W=1u L=180.00n
MM44 net0109 ~D VDD VDD p_18 W=1u L=180.00n
MM43 net0109 ~C VDD VDD p_18 W=1u L=180.00n
MM42 net0109 B VDD VDD p_18 W=1u L=180.00n
MM41 O5 net0111 VDD VDD p_18 W=1u L=180.00n
MM39 net0111 A VDD VDD p_18 W=1u L=180.00n
MM35 net0111 D VDD VDD p_18 W=1u L=180.00n
MM34 net0111 C VDD VDD p_18 W=1u L=180.00n
MM33 net0111 ~B VDD VDD p_18 W=1u L=180.00n
MM32 O6 net067 VDD VDD p_18 W=1u L=180.00n
MM30 net067 A VDD VDD p_18 W=1u L=180.00n
MM26 net067 ~D VDD VDD p_18 W=1u L=180.00n
MM25 net067 C VDD VDD p_18 W=1u L=180.00n
MM24 net067 ~B VDD VDD p_18 W=1u L=180.00n
MM23 O7 net070 VDD VDD p_18 W=1u L=180.00n
MM21 net070 A VDD VDD p_18 W=1u L=180.00n
MM17 net070 D VDD VDD p_18 W=1u L=180.00n
MM16 net070 ~C VDD VDD p_18 W=1u L=180.00n
MM15 net070 ~B VDD VDD p_18 W=1u L=180.00n
MM13 ~D D VDD VDD p_18 W=1u L=180.00n
MM12 ~C C VDD VDD p_18 W=1u L=180.00n
MM10 O8 net18 VDD VDD p_18 W=1u L=180.00n
MM8 ~B B VDD VDD p_18 W=1u L=180.00n
MM6 net18 A VDD VDD p_18 W=1u L=180.00n
MM2 net18 ~D VDD VDD p_18 W=1u L=180.00n
MM1 net18 ~C VDD VDD p_18 W=1u L=180.00n
MM0 net18 ~B VDD VDD p_18 W=1u L=180.00n
MM76 O1 net0143 VSS VSS n_18 W=500.0n L=180.00n
MM74 net0187 D VSS VSS n_18 W=500.0n L=180.00n
MM73 net0188 C net0187 VSS n_18 W=500.0n L=180.00n
MM72 net0143 B net0188 VSS n_18 W=500.0n L=180.00n
MM67 O2 net0145 VSS VSS n_18 W=500.0n L=180.00n
MM65 net0189 ~D VSS VSS n_18 W=500.0n L=180.00n
MM64 net0190 C net0189 VSS n_18 W=500.0n L=180.00n
MM63 net0145 B net0190 VSS n_18 W=500.0n L=180.00n
MM58 O3 net0107 VSS VSS n_18 W=500.0n L=180.00n
MM56 net0191 D VSS VSS n_18 W=500.0n L=180.00n
MM55 net0192 ~C net0191 VSS n_18 W=500.0n L=180.00n
MM54 net0107 B net0192 VSS n_18 W=500.0n L=180.00n
MM49 O4 net0109 VSS VSS n_18 W=500.0n L=180.00n
MM47 net0193 ~D VSS VSS n_18 W=500.0n L=180.00n
MM46 net0194 ~C net0193 VSS n_18 W=500.0n L=180.00n
MM45 net0109 B net0194 VSS n_18 W=500.0n L=180.00n
MM40 O5 net0111 VSS VSS n_18 W=500.0n L=180.00n
MM38 net0195 D VSS VSS n_18 W=500.0n L=180.00n
MM37 net0196 C net0195 VSS n_18 W=500.0n L=180.00n
MM36 net0111 ~B net0196 VSS n_18 W=500.0n L=180.00n
MM31 O6 net067 VSS VSS n_18 W=500.0n L=180.00n
MM29 net0197 ~D VSS VSS n_18 W=500.0n L=180.00n
MM28 net0198 C net0197 VSS n_18 W=500.0n L=180.00n
MM27 net067 ~B net0198 VSS n_18 W=500.0n L=180.00n
MM22 O7 net070 VSS VSS n_18 W=500.0n L=180.00n
MM20 net0199 D VSS VSS n_18 W=500.0n L=180.00n
MM19 net0200 ~C net0199 VSS n_18 W=500.0n L=180.00n
MM18 net070 ~B net0200 VSS n_18 W=500.0n L=180.00n
MM14 ~D D VSS VSS n_18 W=500.0n L=180.00n
MM11 ~C C VSS VSS n_18 W=500.0n L=180.00n
MM9 O8 net18 VSS VSS n_18 W=500.0n L=180.00n
MM7 ~B B VSS VSS n_18 W=500.0n L=180.00n
MM5 net15 ~D VSS VSS n_18 W=500.0n L=180.00n
MM4 net16 ~C net15 VSS n_18 W=500.0n L=180.00n
MM3 net18 ~B net16 VSS n_18 W=500.0n L=180.00n
.ENDS

