.SUBCKT VCO_INV CTRL ~CTRL IN OUT VDD VSS
MM0 netx CTRL VDD VDD p_18 W=14u L=180.00n
MM1 OUT IN netx VDD p_18 W=1u L=180.00n
MM2 OUT IN nety VSS n_18 W=0.5u L=180.00n
MM4 nety ~CTRL VSS VSS n_18 W=5u L=180.00n
.ENDS

.SUBCKT VCO CTRL CTRLB IN VDD VSS
x1 CTRL CTRLB IN net1 VDD VSS VCO_INV
x2 CTRL CTRLB net1 net2 VDD VSS VCO_INV
x3 CTRL CTRLB net2 net3 VDD VSS VCO_INV
x4 CTRL CTRLB net3 net4 VDD VSS VCO_INV
x5 CTRL CTRLB net4 IN VDD VSS VCO_INV
.ENDS

