.SUBCKT NAND6 A B C D E F OUT VDD VSS
MM0 OUT A VDD VDD p_18 W=1.25u L=180.00n
MM1 OUT B VDD VDD p_18 W=1.25u L=180.00n
MM2 OUT C VDD VDD p_18 W=1.25u L=180.00n
MM3 OUT D VDD VDD p_18 W=1.25u L=180.00n
MM4 OUT E VDD VDD p_18 W=1.25u L=180.00n
MM5 OUT F VDD VDD p_18 W=1.25u L=180.00n
MM6 OUT F net4 VSS n_18 W=3.25u L=180.00n
MM7 net4 E net3 VSS n_18 W=3.25u L=180.00n
MM8 net3 D net2 VSS n_18 W=3.25u L=180.00n
MM9 net2 C net1 VSS n_18 W=3.25u L=180.00n
MM10 net1 B net0 VSS n_18 W=3.25u L=180.00n
MM11 net0 A VSS VSS n_18 W=3.25u L=180.00n
.ENDS

.SUBCKT INV IN OUT VDD VSS
MM0 OUT IN VDD VDD p_18 W=20.41u L=180n
MM1 OUT IN VSS VSS n_18 W=10.21u L=180n
.ENDS

.SUBCKT A IN OUT VDD VSS
X1 IN VDD VDD VDD VDD VDD net0 VDD VSS NAND6
X2 net0 OUT VDD VSS INV
.ENDS
