************************************************************************
* auCdl Netlist:
* 
* Library Name:  mylib
* Top Cell Name: PMOS_pass_t
* View Name:     schematic
* Netlisted on:  Apr  3 22:42:46 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: mylib
* Cell Name:    PMOS_pass_t
* View Name:    schematic
************************************************************************

.SUBCKT PMOS_pass_t CLK IN OUT VDD
*.PININFO CLK:I IN:I VDD:I OUT:O
MM0 IN CLK OUT VDD P_18 W=1u L=180.00n
.ENDS

