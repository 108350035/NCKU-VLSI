* File: /home/IC/NCKU/lab1/pb3/decoder.pex.spi
* Created: Mon Apr  7 16:13:16 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.subckt decoder  C A D B O5 O7 O1 O3 O6 O8 VSS VDD O2 O4
* 
MM11 ~C C VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
MM14 ~D D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
MM7 ~B B VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
MM40 O5 NET0111 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
MM22 O7 NET070 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
MM36 NET0111 ~B NET0196 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
MM18 NET070 ~B NET0200 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
MM37 NET0196 C NET0195 VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
MM19 NET0200 ~C NET0199 VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
MM38 NET0195 D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
MM20 NET0199 D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
MM74 NET0187 D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
MM56 NET0191 D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
MM73 NET0188 C NET0187 VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
MM55 NET0192 ~C NET0191 VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
MM72 NET0143 B NET0188 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
MM54 NET0107 B NET0192 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
MM76 O1 NET0143 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
MM58 O3 NET0107 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
MM31 O6 NET067 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
MM9 O8 NET18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
MM27 NET067 ~B NET0198 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
MM3 NET18 ~B NET16 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
MM28 NET0198 C NET0197 VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
MM4 NET16 ~C NET15 VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
MM29 NET0197 ~D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
MM5 NET15 ~D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07
+ PS=1.48e-06
MM65 NET0189 ~D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
MM47 NET0193 ~D VSS VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
MM64 NET0190 C NET0189 VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
MM46 NET0194 ~C NET0193 VSS N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
MM63 NET0145 B NET0190 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
MM45 NET0109 B NET0194 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
MM67 O2 NET0145 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
MM49 O4 NET0109 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
MM12 ~C C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM13 ~D D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM8 ~B B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM41 O5 NET0111 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM23 O7 NET070 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM39 NET0111 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM21 NET070 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM33 NET0111 ~B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13
+ PD=5.1e-07 PS=5.1e-07
MM15 NET070 ~B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM34 NET0111 C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM16 NET070 ~C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM35 NET0111 D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM17 NET070 D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM71 NET0143 D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM53 NET0107 D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM70 NET0143 C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM52 NET0107 ~C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13
+ PD=5.1e-07 PS=5.1e-07
MM69 NET0143 B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM51 NET0107 B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM75 NET0143 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM57 NET0107 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM77 O1 NET0143 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM59 O3 NET0107 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM32 O6 NET067 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM10 O8 NET18 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM30 NET067 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM6 NET18 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM24 NET067 ~B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM0 NET18 ~B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM25 NET067 C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM1 NET18 ~C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM26 NET067 ~D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM2 NET18 ~D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM62 NET0145 ~D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13
+ PD=1.98e-06 PS=5.1e-07
MM44 NET0109 ~D VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13
+ PD=1.98e-06 PS=5.1e-07
MM61 NET0145 C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM43 NET0109 ~C VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13
+ PD=5.1e-07 PS=5.1e-07
MM60 NET0145 B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM42 NET0109 B VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07
+ PS=5.1e-07
MM66 NET0145 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM48 NET0109 A VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
MM68 O2 NET0145 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
MM50 O4 NET0109 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06
+ PS=1.98e-06
c_1 C 0 5.90876f
c_2 A 0 7.87713f
c_3 D 0 3.98888f
c_4 ~B 0 5.78267f
c_5 ~C 0 5.89586f
c_6 ~D 0 4.36898f
c_7 B 0 5.99128f
c_8 O5 0 0.599966f
c_9 O7 0 0.584911f
c_10 NET0111 0 2.22338f
c_11 NET070 0 1.98288f
c_12 NET0143 0 2.12921f
c_13 NET0107 0 2.04791f
c_14 O1 0 0.603073f
c_15 O3 0 0.589041f
c_16 O6 0 0.603084f
c_17 O8 0 0.58904f
c_18 NET067 0 2.19276f
c_19 NET18 0 2.00326f
c_20 NET0145 0 2.01939f
c_21 NET0109 0 1.96709f
c_22 VSS 0 4.3485f
c_23 VDD 0 9.19902f
c_24 O2 0 0.487312f
c_25 O4 0 0.489855f
*
.include "/home/IC/NCKU/lab1/pb3/decoder.pex.spi.DECODER.pxi"
*
.ends
*
*
