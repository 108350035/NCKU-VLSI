************************************************************************
* auCdl Netlist:
* 
* Library Name:  mylib
* Top Cell Name: mux_2to1_2
* View Name:     schematic
* Netlisted on:  Apr  5 21:23:16 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: mylib
* Cell Name:    mux_2to1_2
* View Name:    schematic
************************************************************************

.SUBCKT mux_2to1_2 A0 A1 OUT S VDD VSS
*.PININFO A0:I A1:I S:I VDD:I VSS:I OUT:O
MM10 ~S S VSS VSS n_18 W=500.0n L=180.00n m=1
MM8 OUT net34 VSS VSS n_18 W=500.0n L=180.00n m=1
MM5 net44 A0 VSS VSS n_18 W=500.0n L=180.00n
MM4 net34 ~S net44 VSS n_18 W=500.0n L=180.00n
MM1 net45 A1 VSS VSS n_18 W=500.0n L=180.00n
MM0 net34 S net45 VSS n_18 W=500.0n L=180.00n
MM11 ~S S VDD VDD p_18 W=1u L=180.00n m=1
MM9 OUT net34 VDD VDD p_18 W=1u L=180.00n m=1
MM7 net34 S net43 VDD p_18 W=1u L=180.00n
MM6 net43 A0 VDD VDD p_18 W=1u L=180.00n
MM3 net34 ~S net46 VDD p_18 W=1u L=180.00n
MM2 net46 A1 VDD VDD p_18 W=1u L=180.00n
.ENDS

