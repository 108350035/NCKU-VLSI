.SUBCKT NAND3 A B C OUT VDD VSS
MM0 OUT A VDD VDD p_18 W=2u L=180.00n
MM1 OUT B VDD VDD p_18 W=2u L=180.00n
MM2 OUT C VDD VDD p_18 W=2u L=180.00n
MM3 OUT C net1 VSS n_18 W=3u L=180.00n
MM4 net1 B net0 VSS n_18 W=3u L=180.00n
MM5 net0 A VSS VSS n_18 W=3u L=180.00n
.ENDS

.SUBCKT NAND2 A B OUT VDD VSS
MM0 OUT A VDD VDD p_18 W=22.36u L=180.00n
MM1 OUT B VDD VDD p_18 W=22.36u L=180.00n
MM4 OUT B net0 VSS n_18 W=22.36u L=180.00n
MM5 net0 A VSS VSS n_18 W=22.36u L=180.00n
.ENDS

.SUBCKT INV IN OUT VDD VSS
MM0 OUT IN VDD VDD p_18 W=7.72u L=180n
MM1 OUT IN VSS VSS n_18 W=3.86u L=180n
.ENDS

.SUBCKT INV2 IN OUT VDD VSS
MM0 OUT IN VDD VDD p_18 W=86.3u L=180n
MM1 OUT IN VSS VSS n_18 W=43.1u L=180n
.ENDS

.SUBCKT D IN OUT VDD VSS
X1 VDD VDD VDD net0 VDD VSS NAND3
X2 net0 net1 VDD VSS INV
X3 IN VDD VDD net2 VDD VSS NAND3
X4 net2 net3 VDD VSS INV
X5 net3 net1 net4 VDD VSS NAND2
X6 net4 OUT VDD VSS INV2
.ENDS
