.SUBCKT NOR3 A B C OUT VDD VSS
MM0 net0 A VDD VDD p_18 W=18u L=180.00n
MM1 net1 B net0 VDD p_18 W=18u L=180.00n
MM2 OUT C net1 VDD p_18 W=18u L=180.00n
MM3 OUT C VSS VSS n_18 W=2u L=180.00n
MM4 OUT B VSS VSS n_18 W=2u L=180.00n
MM5 OUT A VSS VSS n_18 W=2u L=180.00n
.ENDS

.SUBCKT NOR3_CHAIN pulse_in pulse_out VDD VSS
X1 VSS VSS pulse_in w0 VDD VSS NOR3
X2 VSS VSS w0 IN VDD VSS NOR3 M=M1
X3 VSS VSS IN OUT VDD VSS NOR3 M=M2
X4 VSS VSS OUT w1 VDD VSS NOR3 M=M3
X5 VSS VSS w1 pulse_out VDD VSS NOR3 M=M4
.ENDS

