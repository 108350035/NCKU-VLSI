* File: AND6_domino.pex.spi
* Created: Tue Apr 22 14:26:13 2025
* Program "Calibre xRC"
* Version "v2019.3_15.11"
* 
.include "AND6_domino.pex.spi.pex"
.subckt nand6  CLK F E D C B A VDD OUT VSS
* 
* VSS	VSS
* OUT	OUT
* VDD	VDD
* A	A
* B	B
* C	C
* D	D
* E	E
* F	F
* CLK	CLK
MM9 N_NETY_MM9_d N_F_MM9_g N_NET5_MM9_s N_VSS_MM9_b N_18 L=1.8e-07 W=2.7e-06
+ AD=1.323e-12 AS=6.75e-13 PD=3.68e-06 PS=5e-07
MM8 N_NET5_MM8_d N_E_MM8_g N_NET4_MM8_s N_VSS_MM9_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.75e-13 AS=6.75e-13 PD=5e-07 PS=5e-07
MM7 N_NET4_MM7_d N_D_MM7_g N_NET3_MM7_s N_VSS_MM9_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.75e-13 AS=6.75e-13 PD=5e-07 PS=5e-07
MM6 N_NET3_MM6_d N_CLK_MM6_g N_VSS_MM6_s N_VSS_MM9_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.75e-13 AS=1.323e-12 PD=5e-07 PS=3.68e-06
MM4 N_NETX_MM4_d N_C_MM4_g N_NET2_MM4_s N_VSS_MM9_b N_18 L=1.8e-07 W=2.7e-06
+ AD=1.323e-12 AS=6.75e-13 PD=3.68e-06 PS=5e-07
MM3 N_NET2_MM3_d N_B_MM3_g N_NET1_MM3_s N_VSS_MM9_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.75e-13 AS=6.75e-13 PD=5e-07 PS=5e-07
MM2 N_NET1_MM2_d N_A_MM2_g N_NET0_MM2_s N_VSS_MM9_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.75e-13 AS=6.75e-13 PD=5e-07 PS=5e-07
MM1 N_NET0_MM1_d N_CLK_MM1_g N_VSS_MM1_s N_VSS_MM9_b N_18 L=1.8e-07 W=2.7e-06
+ AD=6.75e-13 AS=1.323e-12 PD=5e-07 PS=3.68e-06
MM12 N_OUT_MM12_d N_NETX_MM12_g N_VSS_MM12_s N_VSS_MM9_b N_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
MM13 N_OUT_MM13_d N_NETY_MM13_g N_VSS_MM13_s N_VSS_MM9_b N_18 L=1.8e-07 W=1e-06
+ AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
MM5 N_NETY_MM5_d N_CLK_MM5_g N_VDD_MM5_s N_VDD_MM5_b P_18 L=1.8e-07 W=6.8e-07
+ AD=3.332e-13 AS=3.332e-13 PD=1.66e-06 PS=1.66e-06
MM0 N_NETX_MM0_d N_CLK_MM0_g N_VDD_MM0_s N_VDD_MM5_b P_18 L=1.8e-07 W=6.8e-07
+ AD=3.332e-13 AS=3.332e-13 PD=1.66e-06 PS=1.66e-06
MM10 N_NET6_MM10_d N_NETX_MM10_g N_VDD_MM10_s N_VDD_MM5_b P_18 L=1.8e-07 W=2e-06
+ AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07
MM10@4 N_NET6_MM10@4_d N_NETX_MM10@4_g N_VDD_MM10@4_s N_VDD_MM5_b P_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM10@3 N_NET6_MM10@3_d N_NETX_MM10@3_g N_VDD_MM10@3_s N_VDD_MM5_b P_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM10@2 N_NET6_MM10@2_d N_NETX_MM10@2_g N_VDD_MM10@2_s N_VDD_MM5_b P_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM11 N_OUT_MM11_d N_NETY_MM11_g N_NET6_MM11_s N_VDD_MM5_b P_18 L=1.8e-07 W=2e-06
+ AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM11@4 N_OUT_MM11@4_d N_NETY_MM11@4_g N_NET6_MM11@4_s N_VDD_MM5_b P_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM11@3 N_OUT_MM11@3_d N_NETY_MM11@3_g N_NET6_MM11@3_s N_VDD_MM5_b P_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM11@2 N_OUT_MM11@2_d N_NETY_MM11@2_g N_NET6_MM11@2_s N_VDD_MM5_b P_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06
*
.include "AND6_domino.pex.spi.AND6_DOMINO.pxi"
*
.ends
*
*
